module cache_decoder(out[4095:0], line_select[11:0]);
	input [11:0] line_select;
	output [4095:0] out;
endmodule